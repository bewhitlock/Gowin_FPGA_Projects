module dot_clock_gen (
    input board, 
    output dotclock
);
assign dotclock = board;
endmodule